***Include Library****


***create Instance***
*name node1 node2 value*
R1 1 2 1k
R2 2 0 1k
V  1 0 5


***perform operations***

.op
.end

